-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 15.1.1 Build 189 12/02/2015 SJ Lite Edition
-- Created on Tue Apr 18 19:21:32 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DrinksMachineFSM IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        coin20 : IN STD_LOGIC := '0';
        coin50 : IN STD_LOGIC := '0';
        drink : OUT STD_LOGIC
    );
END DrinksMachineFSM;

ARCHITECTURE BEHAVIOR OF DrinksMachineFSM IS
    TYPE type_fstate IS (st0,st1,st2,st3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,coin20,coin50)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= st0;
            drink <= '0';
        ELSE
            drink <= '0';
            CASE fstate IS
                WHEN st0 =>
                    IF (((coin20 = '0') AND (coin50 = '0'))) THEN
                        reg_fstate <= st0;
                    ELSIF (((coin20 = '1') AND (coin50 = '0'))) THEN
                        reg_fstate <= st1;
                    ELSIF ((coin50 = '1')) THEN
                        reg_fstate <= st2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st0;
                    END IF;

                    drink <= '0';
                WHEN st1 =>
                    IF (((coin20 = '0') AND (coin50 = '0'))) THEN
                        reg_fstate <= st1;
                    ELSIF (((coin20 = '1') AND (coin50 = '0'))) THEN
                        reg_fstate <= st2;
                    ELSIF ((coin50 = '1')) THEN
                        reg_fstate <= st3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st1;
                    END IF;

                    drink <= '0';
                WHEN st2 =>
                    IF (((coin20 = '0') AND (coin50 = '0'))) THEN
                        reg_fstate <= st2;
                    ELSIF (((coin20 = '1') OR (coin50 = '1'))) THEN
                        reg_fstate <= st3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= st2;
                    END IF;

                    drink <= '0';
                WHEN st3 =>
                    reg_fstate <= st0;

                    drink <= '1';
                WHEN OTHERS => 
                    drink <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
